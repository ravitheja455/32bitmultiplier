`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:09:49 07/05/2013 
// Design Name: 
// Module Name:    MUL16 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MUL16(a, b, p);
    input [15:0] a;
    input [15:0] b;
    output [31:0] p;
assign p[0]=a[0]&b[0];
VER16 v1(1'b0,1'b0,1'b0,1'b0,(a[1]&b[0]),(a[0]&b[1]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[1],x3,x2,x1,x0);
VER16 v2(x3,x2,x1,x0,(a[2]&b[0]),(a[1]&b[1]),(a[0]&b[2]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, p[2],x7,x6,x5,x4);
VER16 v3(x7,x6,x5,x4,(a[3]&b[0]),(a[2]&b[1]),(a[1]&b[2]),(a[0]&b[3]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[3],x11,x10,x9,x8);
VER16 v4(x11,x10,x9,x8,(a[4]&b[0]),(a[3]&b[1]),(a[2]&b[2]),(a[1]&b[3]),(a[0]&b[4]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[4],x15,x14,x13,x12);
VER16 v5(x15,x14,x13,x12,(a[5]&b[0]),(a[4]&b[1]),(a[3]&b[2]),(a[2]&b[3]),(a[1]&b[4]),(a[0]&b[5]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[5],x19,x18,x17,x16);
VER16 v6(x19,x18,x17,x16,(a[6]&b[0]),(a[5]&b[1]),(a[4]&b[2]),(a[3]&b[3]),(a[2]&b[4]),(a[1]&b[5]),(a[0]&b[6]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[6],x23,x22,x21,x20);
VER16 v7(x23,x22,x21,x20,(a[7]&b[0]),(a[6]&b[1]),(a[5]&b[2]),(a[4]&b[3]),(a[3]&b[4]),(a[2]&b[5]),(a[1]&b[6]),(a[0]&b[7]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[7],x27,x26,x25,x24);
VER16 v8(x27,x26,x25,x24,(a[8]&b[0]),(a[7]&b[1]),(a[6]&b[2]),(a[5]&b[3]),(a[4]&b[4]),(a[3]&b[5]),(a[2]&b[6]),(a[1]&b[7]),(a[0]&b[8]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[8],x31,x30,x29,x28);
VER16 v9(x31,x30,x29,x28,(a[9]&b[0]),(a[8]&b[1]),(a[7]&b[2]),(a[6]&b[3]),(a[5]&b[4]),(a[4]&b[5]),(a[3]&b[6]),(a[2]&b[7]),(a[1]&b[8]),(a[0]&b[9]),1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[9],x35,x34,x33,x32);
VER16 v10(x35,x34,x33,x32,(a[10]&b[0]),(a[9]&b[1]),(a[8]&b[2]),(a[7]&b[3]),(a[6]&b[4]),(a[5]&b[5]),(a[4]&b[6]),(a[3]&b[7]),(a[2]&b[8]),(a[1]&b[9]),(a[0]&b[10]),1'b0,1'b0,1'b0,1'b0,1'b0,p[10],x39,x38,x37,x36);
VER16 v11(x39,x38,x37,x36,(a[11]&b[0]),(a[10]&b[1]),(a[9]&b[2]),(a[8]&b[3]),(a[7]&b[4]),(a[6]&b[5]),(a[5]&b[6]),(a[4]&b[7]),(a[3]&b[8]),(a[2]&b[9]),(a[1]&b[10]),(a[0]&b[11]),1'b0,1'b0,1'b0,1'b0,p[11],x43,x42,x41,x40);
VER16 v12(x43,x42,x41,x40,(a[12]&b[0]),(a[11]&b[1]),(a[10]&b[2]),(a[9]&b[3]),(a[8]&b[4]),(a[7]&b[5]),(a[6]&b[6]),(a[5]&b[7]),(a[4]&b[8]),(a[3]&b[9]),(a[2]&b[10]),(a[1]&b[11]),(a[0]&b[12]),1'b0,1'b0,1'b0,p[12],x47,x46,x45,x44);
VER16 v13(x47,x46,x45,x44,(a[13]&b[0]),(a[12]&b[1]),(a[11]&b[2]),(a[10]&b[3]),(a[9]&b[4]),(a[8]&b[5]),(a[7]&b[6]),(a[6]&b[7]),(a[5]&b[8]),(a[4]&b[9]),(a[3]&b[10]),(a[2]&b[11]),(a[1]&b[12]),(a[0]&b[13]),1'b0,1'b0,p[13],x51,x50,x49,x48);
VER16 v14(x51,x50,x49,x48,(a[14]&b[0]),(a[13]&b[1]),(a[12]&b[2]),(a[11]&b[3]),(a[10]&b[4]),(a[9]&b[5]),(a[8]&b[6]),(a[7]&b[7]),(a[6]&b[8]),(a[5]&b[9]),(a[4]&b[10]),(a[3]&b[11]),(a[2]&b[12]),(a[1]&b[13]),(a[0]&b[14]),1'b0,p[14],x55,x54,x53,x52);
VER16 v15(x55,x54,x53,x52,(a[15]&b[0]),(a[14]&b[1]),(a[13]&b[2]),(a[12]&b[3]),(a[11]&b[4]),(a[10]&b[5]),(a[9]&b[6]),(a[8]&b[7]),(a[7]&b[8]),(a[6]&b[9]),(a[5]&b[10]),(a[4]&b[11]),(a[3]&b[12]),(a[2]&b[13]),(a[1]&b[14]),(a[0]&b[15]),p[15],x59,x58,x57,x56);
VER16 v16(x59,x58,x57,x56,1'b0,(a[15]&b[1]),(a[14]&b[2]),(a[13]&b[3]),(a[12]&b[4]),(a[11]&b[5]),(a[10]&b[6]),(a[9]&b[7]),(a[8]&b[8]),(a[7]&b[9]),(a[6]&b[10]),(a[5]&b[11]),(a[4]&b[12]),(a[3]&b[13]),(a[2]&b[14]),(a[1]&b[15]),p[16],x63,x62,x61,x60);
VER16 v17(x63,x62,x61,x60,1'b0,1'b0,(a[15]&b[2]),(a[14]&b[3]),(a[13]&b[4]),(a[12]&b[5]),(a[11]&b[6]),(a[10]&b[7]),(a[9]&b[8]),(a[8]&b[9]),(a[7]&b[10]),(a[6]&b[11]),(a[5]&b[12]),(a[4]&b[13]),(a[3]&b[14]),(a[2]&b[15]),p[17],x67,x66,x65,x64);
VER16 v18(x67,x66,x65,x64,1'b0,1'b0,1'b0,(a[15]&b[3]),(a[14]&b[4]),(a[13]&b[5]),(a[12]&b[6]),(a[11]&b[7]),(a[10]&b[8]),(a[9]&b[9]),(a[8]&b[10]),(a[7]&b[11]),(a[6]&b[12]),(a[5]&b[13]),(a[4]&b[14]),(a[3]&b[15]),p[18],x71,x70,x69,x68);
VER16 v19(x71,x70,x69,x68,1'b0,1'b0,1'b0,1'b0,(a[15]&b[4]),(a[14]&b[5]),(a[13]&b[6]),(a[12]&b[7]),(a[11]&b[8]),(a[10]&b[9]),(a[9]&b[10]),(a[8]&b[11]),(a[7]&b[12]),(a[6]&b[13]),(a[5]&b[14]),(a[4]&b[15]),p[19],x75,x74,x73,x72);
VER16 v20(x75,x74,x73,x72,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[5]),(a[14]&b[6]),(a[13]&b[7]),(a[12]&b[8]),(a[11]&b[9]),(a[10]&b[10]),(a[9]&b[11]),(a[8]&b[12]),(a[7]&b[13]),(a[6]&b[14]),(a[5]&b[15]),p[20],x79,x78,x77,x76);
VER16 v21(x79,x78,x77,x76,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[6]),(a[14]&b[7]),(a[13]&b[8]),(a[12]&b[9]),(a[11]&b[10]),(a[10]&b[11]),(a[9]&b[12]),(a[8]&b[13]),(a[7]&b[14]),(a[6]&b[15]),p[21],x83,x82,x81,x80);
VER16 v22(x83,x82,x81,x80,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[7]),(a[14]&b[8]),(a[13]&b[9]),(a[12]&b[10]),(a[11]&b[11]),(a[10]&b[12]),(a[9]&b[13]),(a[8]&b[14]),(a[7]&b[15]),p[22],x87,x86,x85,x84);
VER16 v23(x87,x86,x85,x84,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[8]),(a[14]&b[9]),(a[13]&b[10]),(a[12]&b[11]),(a[11]&b[12]),(a[10]&b[13]),(a[9]&b[14]),(a[8]&b[15]),p[23],x91,x90,x89,x88);
VER16 v24(x91,x90,x89,x88,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[9]),(a[14]&b[10]),(a[13]&b[11]),(a[12]&b[12]),(a[11]&b[13]),(a[10]&b[14]),(a[9]&b[15]),p[24],x95,x94,x93,x92);
VER16 v25(x95,x94,x93,x92,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[10]),(a[14]&b[11]),(a[13]&b[12]),(a[12]&b[13]),(a[11]&b[14]),(a[10]&b[15]),p[25],x99,x98,x97,x96);
VER16 v26(x99,x98,x97,x96,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[11]),(a[14]&b[12]),(a[13]&b[13]),(a[12]&b[14]),(a[11]&b[15]),p[26],x103,x102,x101,x100);
VER16 v27(x103,x102,x101,x100,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[12]),(a[14]&b[13]),(a[13]&b[14]),(a[12]&b[15]),p[27],x107,x106,x105,x104);
VER16 v28(x107,x106,x105,x104,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[13]),(a[14]&b[14]),(a[13]&b[15]),p[28],x111,x110,x109,x108);
VER16 v29(x111,x110,x109,x108,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[14]),(a[14]&b[15]),p[29],x115,x114,x113,x112);
VER16 v30(x115,x114,x113,x112,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,(a[15]&b[15]),p[30],x119,x118,x117,x116);
VER16 v31(x119,x118,x117,x116,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,p[31],x123,x122,x121,x120);
endmodule
